library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity memory is
Port ( 
	dir : in STD_LOGIC_VECTOR (11 downto 0);
	data : out STD_LOGIC_VECTOR (97 downto 0));
end memory;

architecture Behavioral of memory is

begin
	process(dir)
	begin
	
		-- DATA FORMAT
		-- |    PRUEBA    |VF| Ins |                LIGA                 |
		--  P4 P3 P2 P1 P0 VF I1 I0 L11 L10 L9 L8 L7 L6 L5 L4 L3 L2 L1 L0 nCRI EB1 EB0 nWB EA1 EA0 nWA selbus UPA9 UPA8 UPA7 UPA6 UPA5 UPA4 UPA3 UPA2 UPA1 UPA0 nOEUPA nDUPA selmux nEX2 nEX1 nEX0 X2 X1 X0 EnaY nERA2 nERA1 nERA0 RA2 RA1 RA0 nEAP2 nEAP1 nEAP0 AP2 AP1 AP0 nEPC2 nEPC1 nEPC0 PC2 PC1 PC0 nCBD nAS nRW BD DINT HINT SET_IRQ SET_XIRQ B9 B8 B7 B6 B5 B4 B3 B2 B1 B0 CC CN CV CZ CI CH CX CS nHB ACCSEC

		-- Cadena por default: "00000" & "0" & "00" & "000000000000" & "10010010000000000011011100001110001110001110001110000000000000000000000010"
		
		--if(dir=    X"000") then data <= "00000" & "0" & "00" & "000000000000" & "10010010000000000011011100001110001110001110001110000000000000000000000010";
		--elsif(dir= X"001") then data <= "00000" & "0" & "00" & "000000000000" & "00000000000000000000000000000000000000000000000000000000000000000000000000"; 

		--INITIALIZATION STATES (000 - 007) HARD CODE
		if(dir=    X"000") then data <= "11000001000000001000100100100000000000110111000011100011100011100011111110000000000000000000000010";

		--FETCH										  
		elsif(dir= X"008") then data <= "00000000000000000000100100100000000000110111000011100011100001100001111110000000000000000000000010";
		elsif(dir= X"009") then data <= "00000000000000000000000100100000000000110111000011100011100011100111111010000000000000000000000010";
		elsif(dir= X"00A") then data <= "00000010000000000000100100100000000000110111000011100011100011100011111110000000000000000000000010";

		--LDAA (INM)
		elsif(dir= X"860") then data <= "00000000000000000000100100100000000000110111000011100011100001100001111110000000000000000000000010";
		elsif(dir= X"861") then data <= "00000000000000000000100101000000000000110111000011100011100011100111111010000000000000000000000010";
		elsif(dir= X"862") then data <= "01111111000000000000100100100000000000110111000011100011100011100011111110000000010011000111000010";
		elsif(dir= X"863") then data <= "11000001000000001001100100100000000000110111000011100011100001100001111110000000000000000000000010";

		--LDAB (INM)
		elsif(dir= X"C60") then data <= "00000000000000000000100100100000000000110111000011100011100001100001111110000000000000000000000010";
		elsif(dir= X"C61") then data <= "00000000000000000000101000100000000000110111000011100011100011100111111010000000000000000000000010";
		elsif(dir= X"C62") then data <= "01111111000000000000100100100000000000110111000011100011100011100011111110000000100101000111000010";
		elsif(dir= X"C63") then data <= "11000001000000001001100100100000000000110111000011100011100001100001111110000000000000000000000010";

		--ABA (INH)
		elsif(dir= X"1B0") then data <= "00000000000000000000111111100000000001111111000011100011100011100011111110000000000000000000000010";
		elsif(dir= X"1B1") then data <= "01111111000000000000100101000000000000000111000011100011100011100011111110000000000000001111010010";
		elsif(dir= X"1B2") then data <= "11000001000000001001100100100000000000110111000011100011100001100001111110000000000000000000000010";

		--JMP (EXT)
		elsif(dir= X"7E0") then data <= "00000000000000000000100100100000000000110111000011100011100001100001111110000000000000000000000010";
		elsif(dir= X"7E1") then data <= "00000000000000000000100100100000000000110111000010110011100011100111111011000000000000000000000010";
		elsif(dir= X"7E2") then data <= "00000000000000000000100100100000000000110111000011100011100001100001111110000000000000000000000010";
		elsif(dir= X"7E3") then data <= "00000000000000000000100100100000000000110111000011001111100011100111111010000000000000000000000010";
		elsif(dir= X"7E4") then data <= "01111111000000000000100100100000000000110111000010000011100010010111111110000000000000000000000010";
		elsif(dir= X"7E5") then data <= "11000001000000001001100100100000000000110111000011100011100001100001111110000000000000000000000010";

		--CMP (INH)
		elsif(dir = X"1A0") then data <= "00000000000000000000111111100000100001111111000011100011100011100011111110000000000000000000000011";
		elsif(dir = X"1A1") then data <= "01111111000000000000100100100000000000000111000011100011100011100011111110000000000000001111010010";
		elsif(dir = X"1A2") then data <= "11000001000000001001100100100000000000110111000011100011100001100001111110000000000000000000000010";

		--JE (EXT)
		elsif(dir = X"7D0") then data <= "00000000000000000000100100100000000000110111000011100011100001100001111110000000000000000000000010";
		elsif(dir = X"7D1") then data <= "00000000000000000000100100100000000000110111000010110011100011100111111011000000000000000000000010";
		elsif(dir = X"7D2") then data <= "00000000000000000000100100100000000000110111000011100011100001100001111110000000000000000000000010";
		elsif(dir = X"7D3") then data <= "10010001011111010101100100100000000000110111000011001111100011100111111010000000000000000000000010";
		elsif(dir = X"7D4") then data <= "01111111000000000000100100100000000000110111000010000011100010010111111110000000000000000000000010";
		elsif(dir = X"7D5") then data <= "11000001000000000000100100100000000000110111000011100011100001100001111110000000000000000000000010";

		--LDX (INS)
		elsif(dir = X"5B0") then data <= "00000000000000000000100100100000000000110111000011100011100001100001111110000000000000000000000010";
		elsif(dir = X"5B1") then data <= "00000000000000000000100100100000000000110101100011100011100011100111111110000000000000000000000010";
		elsif(dir = X"5B2") then data <= "00000000000000000000100100100000000000110111000011100011100001100001111110000000000000000000000010";
		
		elsif(dir = X"5B3") then data <= "00000000000000000000100100100000000000110110011011100011100011100111111110000000000000000000000010";
		elsif(dir = X"5B4") then data <= "01111111000000000000100100100000000000110111000011100011100011100011111110000000110111000111000010";
		elsif(dir = X"5B5") then data <= "11000001000000001001100100100000000000110111000011100011100001100001111110000000000000000000000010";

		--LDAA (DIR)
		elsif(dir = X"A90") then data <= "00000000000000000000100111100001000000110111000011100011100011100011111110000000000000000000000010";
		elsif(dir = X"A91") then data <= "00000000000000000000100100100000000000000111000010110011100011100011111110000000000000000000000010";
		elsif(dir = X"A92") then data <= "00000000000000000000100100100000000000110111000011100011100001100001111110000000000000000000000010";
		elsif(dir = X"A93") then data <= "00000000000000000000100100100000000000110111000011001111100011100111111010000000000000000000000010";
		elsif(dir = X"A94") then data <= "00000000000000000000100100100000000000110111000001100011100011100001111110000000000000000000000010";
		elsif(dir = X"A95") then data <= "00000000000000000000100101000000000000110111000011100011100011100111111010000000000000000000000010";
		elsif(dir = X"A96") then data <= "01111111000000000000100100100000000000110111000011100011100011100011111110000000010011000111000010";
		elsif(dir = X"A97") then data <= "11000001000000001001100100100000000000110111000011100011100001100001111110000000000000000000000010";

		--LDAB (DIR)
		elsif(dir = X"AA0") then data <= "00000000000000000000100111100001000000110111000011100011100011100011111110000000000000000000000010";
		elsif(dir = X"AA1") then data <= "00000000000000000000100100100000000000000111000010110011100011100011111110000000000000000000000010";
		elsif(dir = X"AA2") then data <= "00000000000000000000100100100000000000110111000011100011100001100001111110000000000000000000000010";
		elsif(dir = X"AA3") then data <= "00000000000000000000100100100000000000110111000011001111100011100111111010000000000000000000000010";
		elsif(dir = X"AA4") then data <= "00000000000000000000100100100000000000110111000001100011100011100001111110000000000000000000000010";
		elsif(dir = X"AA5") then data <= "00000000000000000000101000100000000000110111000011100011100011100111111010000000000000000000000010";
		elsif(dir = X"AA6") then data <= "01111111000000000000100100100000000000110111000011100011100011100011111110000000100101000111000010";
		elsif(dir = X"AA7") then data <= "11000001000000001001100100100000000000110111000011100011100001100001111110000000000000000000000010";


		--STAA (DIR)
		elsif(dir = X"A80") then data <= "00000000000000000000100111100001000000110111000011100011100011100011111110000000000000000000000010";
		elsif(dir = X"A81") then data <= "00000000000000000000100100100000000000000111000010110011100011100011111110000000000000000000000010";
		elsif(dir = X"A82") then data <= "00000000000000000000100100100000000000110111000011100011100001100001111110000000000000000000000010";
		elsif(dir = X"A83") then data <= "00000000000000000000100100100000000000110111000011001111100011100111111010000000000000000000000010";
		elsif(dir = X"A84") then data <= "00000000000000000000100100100000000000110111000001100011100011100001111110000000000000000000000010";
		elsif(dir = X"A85") then data <= "00000000000000000000100101100000000000110111000011100011100011100011111000000000000000000000000010";
		elsif(dir = X"A86") then data <= "01111111000000000000100100100000000000110111000011100011100011100011111110000000010011000111000010";
		elsif(dir = X"A87") then data <= "11000001000000001001100100100000000000110111000011100011100001100001111110000000000000000000000010";

		--STAB (DIR)
		elsif(dir = X"A90") then data <= "00000000000000000000100111100001000000110111000011100011100011100011111110000000000000000000000010";
		elsif(dir = X"A91") then data <= "00000000000000000000100100100000000000000111000010110011100011100011111110000000000000000000000010";
		elsif(dir = X"A92") then data <= "00000000000000000000100100100000000000110111000011100011100001100001111110000000000000000000000010";
		elsif(dir = X"A93") then data <= "00000000000000000000100100100000000000110111000011001111100011100111111010000000000000000000000010";
		elsif(dir = X"A94") then data <= "00000000000000000000100100100000000000110111000001100011100011100001111110000000000000000000000010";
		elsif(dir = X"A95") then data <= "00000000000000000000101100100000000000110111000011100011100011100011111000000000000000000000000010";
		elsif(dir = X"A96") then data <= "01111111000000000000100100100000000000110111000011100011100011100011111110000000100101000111000010";
		elsif(dir = X"A97") then data <= "11000001000000001001100100100000000000110111000011100011100001100001111110000000000000000000000010";


		--ANDA (INM)
		elsif(dir = X"D70") then data <= "00000000000000000000100111100000000000110111000011100011100001100001111110000000000000000000000010";
		elsif(dir = X"D71") then data <= "00000000000000000000100111100101000101110111000011100011100011100111111010000000000000000000000010";
		elsif(dir = X"D72") then data <= "01111111000000000000100100101001000000110111000011100011100011100011111111111100000000000111000010";
		elsif(dir = X"D73") then data <= "11000001000000001001100100100000000000110111000011100011100001100001111110000000000000000000000010";

		--BRA (REL)
		elsif(dir = X"B10") then data <= "00000000000000000000100100100000000000110111000011001111100001100001111110000000000000000000000000";
		elsif(dir = X"B11") then data <= "00000000000000000000100100100000110111110111000011100011100011100111111010000000000000000000000010";
		elsif(dir = X"B12") then data <= "00000000000000000000100100100010000110111111000011100011100011000011111110000000000000000000000010";
		elsif(dir = X"B13") then data <= "00000101000000001000100100100000000000000111000011100011100011001111111110000000000000001000000010";
		elsif(dir = X"B14") then data <= "00000000000000000000100100110010000111110111000011100011100010100011111110000000000000000000000010";
		elsif(dir = X"B15") then data <= "00000000000000000000100100100000000000000111000011100011100010110011111110000000000000000000000010";
		elsif(dir = X"B16") then data <= "01111111000000000000100100100000000000110111000011000011100011100011111110000000000000011000000000";
		elsif(dir = X"B17") then data <= "11000001000000001001100100100000000000110111000011100011100001100001111110000000000000000000000010";
		elsif(dir = X"B18") then data <= "11000001000000000101100100110010100111110111000011100011100010100011111110000000000000000000000010";

		--INCX (INH)
		elsif(dir = X"80") then data <= "00000000000000000000100100100000000000110111001011100011100011100011111110000000000000000000000010";
		elsif(dir = X"81") then data <= "01111111000000000000100100100000000000110111000011100011100011100011111110000000000110000001000010";
		elsif(dir = X"82") then data <= "11000001000000001001100100100000000000110111000011100011100001100001111110000000000000000000000010";

		-- NOP
		elsif(dir = X"10") then data <= "01111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
		elsif(dir = X"11") then data <= "11000001000000001001100100100000000000110111000011100011100001100001111110000000000000000000000010";



		else data <= "00000000000000000000100100100000000000110111000011100011100011100011111110000000000000000000000010";

		end if;
	end process;
end Behavioral;

-- elsif(dir = X"A") then data <= "";